magic
tech sky130A
magscale 1 2
timestamp 1768494946
<< locali >>
rect 213 1960 448 2040
rect -96 -200 96 152
rect 1056 -200 1248 152
rect -200 -211 1400 -200
rect -200 -391 294 -211
rect 474 -391 1400 -211
rect -200 -400 1400 -391
<< viali >>
rect 294 -391 474 -211
<< metal1 >>
rect 160 40 224 3951
rect 672 3694 1157 3886
rect 288 -205 480 3530
rect 965 3078 1157 3694
rect 672 2886 1157 3078
rect 965 1441 1157 2886
rect 672 1249 1158 1441
rect 965 670 1157 1249
rect 676 478 1157 670
rect 672 40 864 120
rect 282 -211 486 -205
rect 282 -391 294 -211
rect 474 -391 486 -211
rect 282 -397 486 -391
use JNWATR_NCH_4C5F0  xo0<0> ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 0
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo0<1>
timestamp 1740610800
transform 1 0 0 0 1 800
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1<0>
timestamp 1740610800
transform 1 0 0 0 1 2400
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1<1>
timestamp 1740610800
transform 1 0 0 0 1 3200
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1
timestamp 1740610800
transform 1 0 0 0 1 1600
box -184 -128 1336 928
<< labels >>
flabel metal1 s 672 40 864 120 0 FreeSans 400 0 0 0 IBNS_20U
port 1 nsew signal bidirectional
flabel metal1 s 288 600 480 680 0 FreeSans 400 0 0 0 VSS
port 2 nsew ground bidirectional
flabel metal1 s 160 360 224 440 0 FreeSans 400 0 0 0 IBPS_5U
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 4000
<< end >>
